type gui_ele_btn_type is array (0 to 29, 0 to 119) of std_logic_vector(11 downto 0);
constant BTN_toggle : gui_ele_btn_type := (
    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"4A1", x"4A1", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"3D1", x"4A1", x"4A1", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"3D1", x"3D1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"4A1", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"4A1", x"4A1", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"4A1", x"4A1", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"4A1", x"4A1", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"4A1", x"4A1", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"070", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF")
);
