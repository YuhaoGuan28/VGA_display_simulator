type gui_ele_font30_type is array (0 to 25, 0 to 19) of std_logic_vector(11 downto 0);
constant A_30 : gui_ele_font30_type := (
    (x"000", x"000", x"000", x"AA0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"AA0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"AA0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"440", x"660", x"880", x"880", x"880", x"880", x"880", x"880", x"880", x"880", x"880", x"330", x"000", x"000", x"000", x"000", x"000"),
    (x"FF0", x"FF0", x"FF0", x"550", x"000", x"220", x"330", x"330", x"330", x"330", x"330", x"330", x"330", x"770", x"FF0", x"FF0", x"FF0", x"000", x"000", x"000"),
    (x"FF0", x"FF0", x"FF0", x"550", x"000", x"110", x"110", x"110", x"110", x"110", x"110", x"110", x"110", x"660", x"FF0", x"FF0", x"FF0", x"000", x"000", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"BB0", x"880", x"880", x"880", x"880", x"880", x"880", x"880", x"880", x"880", x"BB0", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"330", x"330", x"330", x"330", x"330", x"330", x"330", x"330", x"770", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"220", x"110", x"110", x"110", x"110", x"110", x"110", x"110", x"660", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"550", x"FF0", x"FF0", x"FF0", x"330", x"330", x"000"),
    (x"000", x"000", x"330", x"330", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"110", x"330", x"330", x"330", x"000"),
    (x"000", x"000", x"330", x"330", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"110", x"330", x"330", x"330", x"000")
);
