type gui_ele_type is array (0 to 10, 0 to 7) of std_logic_vector(11 downto 0);
    constant Y_12 : gui_ele_font12_type := (
        (x"FF0", x"110", x"000", x"000", x"000", x"FF0", x"110", x"000"),
        (x"770", x"550", x"000", x"000", x"110", x"660", x"440", x"000"),
        (x"000", x"EE0", x"110", x"000", x"FF0", x"110", x"110", x"000"),
        (x"000", x"000", x"660", x"FF0", x"110", x"330", x"000", x"000"),
        (x"000", x"000", x"440", x"FF0", x"440", x"000", x"000", x"000"),
        (x"000", x"000", x"440", x"FF0", x"440", x"000", x"000", x"000"),
        (x"000", x"000", x"440", x"FF0", x"440", x"000", x"000", x"000"),
        (x"000", x"000", x"440", x"FF0", x"440", x"000", x"000", x"000"),
        (x"000", x"000", x"440", x"FF0", x"440", x"000", x"000", x"000"),
        (x"000", x"000", x"440", x"FF0", x"440", x"000", x"000", x"000"),
        (x"000", x"000", x"000", x"110", x"330", x"000", x"000", x"000")
    );
