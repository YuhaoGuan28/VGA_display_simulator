type gui_ele_type is array (0 to 10, 0 to 7) of std_logic_vector(11 downto 0);
    constant J_12 : gui_ele_font12_type := (
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
        (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00")
    );
