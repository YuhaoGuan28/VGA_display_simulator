type gui_ele_type is array (0 to 10, 0 to 7) of std_logic_vector(11 downto 0);
    constant S_12 : gui_ele_font12_type := (
        (x"000", x"EE0", x"FF0", x"FF0", x"FF0", x"FF0", x"110", x"000"),
        (x"110", x"660", x"880", x"880", x"880", x"880", x"440", x"000"),
        (x"FF0", x"110", x"110", x"110", x"110", x"110", x"110", x"000"),
        (x"110", x"FF0", x"FF0", x"FF0", x"FF0", x"000", x"000", x"000"),
        (x"000", x"550", x"880", x"880", x"880", x"CC0", x"000", x"000"),
        (x"000", x"000", x"110", x"110", x"110", x"FF0", x"330", x"000"),
        (x"110", x"000", x"000", x"000", x"000", x"FF0", x"440", x"000"),
        (x"FF0", x"110", x"000", x"000", x"000", x"FF0", x"440", x"000"),
        (x"550", x"880", x"660", x"660", x"660", x"440", x"440", x"000"),
        (x"000", x"EE0", x"FF0", x"FF0", x"FF0", x"110", x"110", x"000"),
        (x"000", x"000", x"330", x"330", x"330", x"330", x"000", x"000")
    );
