type gui_ele_btn_type is array (0 to 29, 0 to 119) of std_logic_vector(11 downto 0);
constant BTN_normal : gui_ele_btn_type := (
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"888", x"888", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"888", x"888", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"FFF", x"FFF", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"888", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"888", x"888", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"888", x"888", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"888", x"888", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"888", x"888", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"555", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000")
);
