type gui_ele_type is array (0 to 25, 0 to 19) of std_logic_vector(11 downto 0);
constant colon_30 : gui_ele_font30_type := (
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"FF0", x"FF0", x"FF0", x"550", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"FF0", x"FF0", x"FF0", x"550", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"660", x"660", x"880", x"550", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"330", x"330", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"110", x"110", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"660", x"660", x"660", x"220", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"FF0", x"FF0", x"FF0", x"550", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"FF0", x"FF0", x"FF0", x"660", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"FF0", x"FF0", x"FF0", x"770", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"330", x"330", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"330", x"330", x"330", x"110", x"000", x"000", x"000", x"000", x"000", x"000", x"000")
);
